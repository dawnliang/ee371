// nios2.v

// Generated using ACDS version 16.0 211

`timescale 1 ps / 1 ps
module nios2 (
		input  wire       clk_clk,                //             clk.clk
		output wire [1:0] ctrl_scanner_export,    //    ctrl_scanner.export
		output wire [1:0] ctrl_sps_export,        //        ctrl_sps.export
		input  wire [1:0] framing_sps_export,     //     framing_sps.export
		input  wire [7:0] in_scanner_export,      //      in_scanner.export
		input  wire [7:0] in_sps_export,          //          in_sps.export
		output wire [7:0] out_scanner_export,     //     out_scanner.export
		output wire [7:0] out_sps_export,         //         out_sps.export
		input  wire       readytotransfer_export, // readytotransfer.export
		input  wire       reset_reset_n           //           reset.reset_n
	);

	wire  [31:0] nios2_qsys_0_data_master_readdata;                            // mm_interconnect_0:nios2_qsys_0_data_master_readdata -> nios2_qsys_0:d_readdata
	wire         nios2_qsys_0_data_master_waitrequest;                         // mm_interconnect_0:nios2_qsys_0_data_master_waitrequest -> nios2_qsys_0:d_waitrequest
	wire         nios2_qsys_0_data_master_debugaccess;                         // nios2_qsys_0:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:nios2_qsys_0_data_master_debugaccess
	wire  [14:0] nios2_qsys_0_data_master_address;                             // nios2_qsys_0:d_address -> mm_interconnect_0:nios2_qsys_0_data_master_address
	wire   [3:0] nios2_qsys_0_data_master_byteenable;                          // nios2_qsys_0:d_byteenable -> mm_interconnect_0:nios2_qsys_0_data_master_byteenable
	wire         nios2_qsys_0_data_master_read;                                // nios2_qsys_0:d_read -> mm_interconnect_0:nios2_qsys_0_data_master_read
	wire         nios2_qsys_0_data_master_write;                               // nios2_qsys_0:d_write -> mm_interconnect_0:nios2_qsys_0_data_master_write
	wire  [31:0] nios2_qsys_0_data_master_writedata;                           // nios2_qsys_0:d_writedata -> mm_interconnect_0:nios2_qsys_0_data_master_writedata
	wire  [31:0] nios2_qsys_0_instruction_master_readdata;                     // mm_interconnect_0:nios2_qsys_0_instruction_master_readdata -> nios2_qsys_0:i_readdata
	wire         nios2_qsys_0_instruction_master_waitrequest;                  // mm_interconnect_0:nios2_qsys_0_instruction_master_waitrequest -> nios2_qsys_0:i_waitrequest
	wire  [14:0] nios2_qsys_0_instruction_master_address;                      // nios2_qsys_0:i_address -> mm_interconnect_0:nios2_qsys_0_instruction_master_address
	wire         nios2_qsys_0_instruction_master_read;                         // nios2_qsys_0:i_read -> mm_interconnect_0:nios2_qsys_0_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;     // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest;  // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;      // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;         // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;    // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata;    // nios2_qsys_0:jtag_debug_module_readdata -> mm_interconnect_0:nios2_qsys_0_jtag_debug_module_readdata
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest; // nios2_qsys_0:jtag_debug_module_waitrequest -> mm_interconnect_0:nios2_qsys_0_jtag_debug_module_waitrequest
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess; // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_debugaccess -> nios2_qsys_0:jtag_debug_module_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address;     // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_address -> nios2_qsys_0:jtag_debug_module_address
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read;        // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_read -> nios2_qsys_0:jtag_debug_module_read
	wire   [3:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable;  // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_byteenable -> nios2_qsys_0:jtag_debug_module_byteenable
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write;       // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_write -> nios2_qsys_0:jtag_debug_module_write
	wire  [31:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata;   // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_writedata -> nios2_qsys_0:jtag_debug_module_writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;             // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;               // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire  [10:0] mm_interconnect_0_onchip_memory2_0_s1_address;                // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;             // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                  // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;              // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                  // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire  [31:0] mm_interconnect_0_in_sps_s1_readdata;                         // in_SPS:readdata -> mm_interconnect_0:in_SPS_s1_readdata
	wire   [1:0] mm_interconnect_0_in_sps_s1_address;                          // mm_interconnect_0:in_SPS_s1_address -> in_SPS:address
	wire         mm_interconnect_0_out_sps_s1_chipselect;                      // mm_interconnect_0:out_SPS_s1_chipselect -> out_SPS:chipselect
	wire  [31:0] mm_interconnect_0_out_sps_s1_readdata;                        // out_SPS:readdata -> mm_interconnect_0:out_SPS_s1_readdata
	wire   [1:0] mm_interconnect_0_out_sps_s1_address;                         // mm_interconnect_0:out_SPS_s1_address -> out_SPS:address
	wire         mm_interconnect_0_out_sps_s1_write;                           // mm_interconnect_0:out_SPS_s1_write -> out_SPS:write_n
	wire  [31:0] mm_interconnect_0_out_sps_s1_writedata;                       // mm_interconnect_0:out_SPS_s1_writedata -> out_SPS:writedata
	wire         mm_interconnect_0_out_scanner_s1_chipselect;                  // mm_interconnect_0:out_scanner_s1_chipselect -> out_scanner:chipselect
	wire  [31:0] mm_interconnect_0_out_scanner_s1_readdata;                    // out_scanner:readdata -> mm_interconnect_0:out_scanner_s1_readdata
	wire   [1:0] mm_interconnect_0_out_scanner_s1_address;                     // mm_interconnect_0:out_scanner_s1_address -> out_scanner:address
	wire         mm_interconnect_0_out_scanner_s1_write;                       // mm_interconnect_0:out_scanner_s1_write -> out_scanner:write_n
	wire  [31:0] mm_interconnect_0_out_scanner_s1_writedata;                   // mm_interconnect_0:out_scanner_s1_writedata -> out_scanner:writedata
	wire  [31:0] mm_interconnect_0_in_scanner_s1_readdata;                     // in_scanner:readdata -> mm_interconnect_0:in_scanner_s1_readdata
	wire   [1:0] mm_interconnect_0_in_scanner_s1_address;                      // mm_interconnect_0:in_scanner_s1_address -> in_scanner:address
	wire         mm_interconnect_0_ctrl_scanner_s1_chipselect;                 // mm_interconnect_0:ctrl_scanner_s1_chipselect -> ctrl_scanner:chipselect
	wire  [31:0] mm_interconnect_0_ctrl_scanner_s1_readdata;                   // ctrl_scanner:readdata -> mm_interconnect_0:ctrl_scanner_s1_readdata
	wire   [1:0] mm_interconnect_0_ctrl_scanner_s1_address;                    // mm_interconnect_0:ctrl_scanner_s1_address -> ctrl_scanner:address
	wire         mm_interconnect_0_ctrl_scanner_s1_write;                      // mm_interconnect_0:ctrl_scanner_s1_write -> ctrl_scanner:write_n
	wire  [31:0] mm_interconnect_0_ctrl_scanner_s1_writedata;                  // mm_interconnect_0:ctrl_scanner_s1_writedata -> ctrl_scanner:writedata
	wire  [31:0] mm_interconnect_0_readytotransfer_s1_readdata;                // readyToTransfer:readdata -> mm_interconnect_0:readyToTransfer_s1_readdata
	wire   [1:0] mm_interconnect_0_readytotransfer_s1_address;                 // mm_interconnect_0:readyToTransfer_s1_address -> readyToTransfer:address
	wire         mm_interconnect_0_ctrl_sps_s1_chipselect;                     // mm_interconnect_0:ctrl_SPS_s1_chipselect -> ctrl_SPS:chipselect
	wire  [31:0] mm_interconnect_0_ctrl_sps_s1_readdata;                       // ctrl_SPS:readdata -> mm_interconnect_0:ctrl_SPS_s1_readdata
	wire   [1:0] mm_interconnect_0_ctrl_sps_s1_address;                        // mm_interconnect_0:ctrl_SPS_s1_address -> ctrl_SPS:address
	wire         mm_interconnect_0_ctrl_sps_s1_write;                          // mm_interconnect_0:ctrl_SPS_s1_write -> ctrl_SPS:write_n
	wire  [31:0] mm_interconnect_0_ctrl_sps_s1_writedata;                      // mm_interconnect_0:ctrl_SPS_s1_writedata -> ctrl_SPS:writedata
	wire  [31:0] mm_interconnect_0_framing_sps_s1_readdata;                    // framing_SPS:readdata -> mm_interconnect_0:framing_SPS_s1_readdata
	wire   [1:0] mm_interconnect_0_framing_sps_s1_address;                     // mm_interconnect_0:framing_SPS_s1_address -> framing_SPS:address
	wire         irq_mapper_receiver0_irq;                                     // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios2_qsys_0_d_irq_irq;                                       // irq_mapper:sender_irq -> nios2_qsys_0:d_irq
	wire         rst_controller_reset_out_reset;                               // rst_controller:reset_out -> [ctrl_SPS:reset_n, ctrl_scanner:reset_n, framing_SPS:reset_n, in_SPS:reset_n, in_scanner:reset_n, irq_mapper:reset, jtag_uart_0:rst_n, mm_interconnect_0:nios2_qsys_0_reset_n_reset_bridge_in_reset_reset, nios2_qsys_0:reset_n, onchip_memory2_0:reset, out_SPS:reset_n, out_scanner:reset_n, readyToTransfer:reset_n, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                           // rst_controller:reset_req -> [nios2_qsys_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	wire         nios2_qsys_0_jtag_debug_module_reset_reset;                   // nios2_qsys_0:jtag_debug_module_resetrequest -> rst_controller:reset_in1

	nios2_ctrl_SPS ctrl_sps (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_ctrl_sps_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_ctrl_sps_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_ctrl_sps_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_ctrl_sps_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_ctrl_sps_s1_readdata),   //                    .readdata
		.out_port   (ctrl_sps_export)                           // external_connection.export
	);

	nios2_ctrl_SPS ctrl_scanner (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_ctrl_scanner_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_ctrl_scanner_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_ctrl_scanner_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_ctrl_scanner_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_ctrl_scanner_s1_readdata),   //                    .readdata
		.out_port   (ctrl_scanner_export)                           // external_connection.export
	);

	nios2_framing_SPS framing_sps (
		.clk      (clk_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_0_framing_sps_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_framing_sps_s1_readdata), //                    .readdata
		.in_port  (framing_sps_export)                         // external_connection.export
	);

	nios2_in_SPS in_sps (
		.clk      (clk_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_0_in_sps_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_in_sps_s1_readdata), //                    .readdata
		.in_port  (in_sps_export)                         // external_connection.export
	);

	nios2_in_SPS in_scanner (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_0_in_scanner_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_in_scanner_s1_readdata), //                    .readdata
		.in_port  (in_scanner_export)                         // external_connection.export
	);

	nios2_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	nios2_nios2_qsys_0 nios2_qsys_0 (
		.clk                                   (clk_clk),                                                      //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                              //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                           //                          .reset_req
		.d_address                             (nios2_qsys_0_data_master_address),                             //               data_master.address
		.d_byteenable                          (nios2_qsys_0_data_master_byteenable),                          //                          .byteenable
		.d_read                                (nios2_qsys_0_data_master_read),                                //                          .read
		.d_readdata                            (nios2_qsys_0_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (nios2_qsys_0_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (nios2_qsys_0_data_master_write),                               //                          .write
		.d_writedata                           (nios2_qsys_0_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (nios2_qsys_0_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (nios2_qsys_0_instruction_master_address),                      //        instruction_master.address
		.i_read                                (nios2_qsys_0_instruction_master_read),                         //                          .read
		.i_readdata                            (nios2_qsys_0_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (nios2_qsys_0_instruction_master_waitrequest),                  //                          .waitrequest
		.d_irq                                 (nios2_qsys_0_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_qsys_0_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                              // custom_instruction_master.readra
	);

	nios2_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)                //       .reset_req
	);

	nios2_out_SPS out_sps (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_out_sps_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_out_sps_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_out_sps_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_out_sps_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_out_sps_s1_readdata),   //                    .readdata
		.out_port   (out_sps_export)                           // external_connection.export
	);

	nios2_out_SPS out_scanner (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_out_scanner_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_out_scanner_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_out_scanner_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_out_scanner_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_out_scanner_s1_readdata),   //                    .readdata
		.out_port   (out_scanner_export)                           // external_connection.export
	);

	nios2_readyToTransfer readytotransfer (
		.clk      (clk_clk),                                       //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address  (mm_interconnect_0_readytotransfer_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_readytotransfer_s1_readdata), //                    .readdata
		.in_port  (readytotransfer_export)                         // external_connection.export
	);

	nios2_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                    (clk_clk),                                                      //                                  clk_0_clk.clk
		.nios2_qsys_0_reset_n_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                               // nios2_qsys_0_reset_n_reset_bridge_in_reset.reset
		.nios2_qsys_0_data_master_address                 (nios2_qsys_0_data_master_address),                             //                   nios2_qsys_0_data_master.address
		.nios2_qsys_0_data_master_waitrequest             (nios2_qsys_0_data_master_waitrequest),                         //                                           .waitrequest
		.nios2_qsys_0_data_master_byteenable              (nios2_qsys_0_data_master_byteenable),                          //                                           .byteenable
		.nios2_qsys_0_data_master_read                    (nios2_qsys_0_data_master_read),                                //                                           .read
		.nios2_qsys_0_data_master_readdata                (nios2_qsys_0_data_master_readdata),                            //                                           .readdata
		.nios2_qsys_0_data_master_write                   (nios2_qsys_0_data_master_write),                               //                                           .write
		.nios2_qsys_0_data_master_writedata               (nios2_qsys_0_data_master_writedata),                           //                                           .writedata
		.nios2_qsys_0_data_master_debugaccess             (nios2_qsys_0_data_master_debugaccess),                         //                                           .debugaccess
		.nios2_qsys_0_instruction_master_address          (nios2_qsys_0_instruction_master_address),                      //            nios2_qsys_0_instruction_master.address
		.nios2_qsys_0_instruction_master_waitrequest      (nios2_qsys_0_instruction_master_waitrequest),                  //                                           .waitrequest
		.nios2_qsys_0_instruction_master_read             (nios2_qsys_0_instruction_master_read),                         //                                           .read
		.nios2_qsys_0_instruction_master_readdata         (nios2_qsys_0_instruction_master_readdata),                     //                                           .readdata
		.ctrl_scanner_s1_address                          (mm_interconnect_0_ctrl_scanner_s1_address),                    //                            ctrl_scanner_s1.address
		.ctrl_scanner_s1_write                            (mm_interconnect_0_ctrl_scanner_s1_write),                      //                                           .write
		.ctrl_scanner_s1_readdata                         (mm_interconnect_0_ctrl_scanner_s1_readdata),                   //                                           .readdata
		.ctrl_scanner_s1_writedata                        (mm_interconnect_0_ctrl_scanner_s1_writedata),                  //                                           .writedata
		.ctrl_scanner_s1_chipselect                       (mm_interconnect_0_ctrl_scanner_s1_chipselect),                 //                                           .chipselect
		.ctrl_SPS_s1_address                              (mm_interconnect_0_ctrl_sps_s1_address),                        //                                ctrl_SPS_s1.address
		.ctrl_SPS_s1_write                                (mm_interconnect_0_ctrl_sps_s1_write),                          //                                           .write
		.ctrl_SPS_s1_readdata                             (mm_interconnect_0_ctrl_sps_s1_readdata),                       //                                           .readdata
		.ctrl_SPS_s1_writedata                            (mm_interconnect_0_ctrl_sps_s1_writedata),                      //                                           .writedata
		.ctrl_SPS_s1_chipselect                           (mm_interconnect_0_ctrl_sps_s1_chipselect),                     //                                           .chipselect
		.framing_SPS_s1_address                           (mm_interconnect_0_framing_sps_s1_address),                     //                             framing_SPS_s1.address
		.framing_SPS_s1_readdata                          (mm_interconnect_0_framing_sps_s1_readdata),                    //                                           .readdata
		.in_scanner_s1_address                            (mm_interconnect_0_in_scanner_s1_address),                      //                              in_scanner_s1.address
		.in_scanner_s1_readdata                           (mm_interconnect_0_in_scanner_s1_readdata),                     //                                           .readdata
		.in_SPS_s1_address                                (mm_interconnect_0_in_sps_s1_address),                          //                                  in_SPS_s1.address
		.in_SPS_s1_readdata                               (mm_interconnect_0_in_sps_s1_readdata),                         //                                           .readdata
		.jtag_uart_0_avalon_jtag_slave_address            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),      //              jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write              (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),        //                                           .write
		.jtag_uart_0_avalon_jtag_slave_read               (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),         //                                           .read
		.jtag_uart_0_avalon_jtag_slave_readdata           (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),     //                                           .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),    //                                           .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest),  //                                           .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),   //                                           .chipselect
		.nios2_qsys_0_jtag_debug_module_address           (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address),     //             nios2_qsys_0_jtag_debug_module.address
		.nios2_qsys_0_jtag_debug_module_write             (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write),       //                                           .write
		.nios2_qsys_0_jtag_debug_module_read              (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read),        //                                           .read
		.nios2_qsys_0_jtag_debug_module_readdata          (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata),    //                                           .readdata
		.nios2_qsys_0_jtag_debug_module_writedata         (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata),   //                                           .writedata
		.nios2_qsys_0_jtag_debug_module_byteenable        (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable),  //                                           .byteenable
		.nios2_qsys_0_jtag_debug_module_waitrequest       (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest), //                                           .waitrequest
		.nios2_qsys_0_jtag_debug_module_debugaccess       (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess), //                                           .debugaccess
		.onchip_memory2_0_s1_address                      (mm_interconnect_0_onchip_memory2_0_s1_address),                //                        onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                        (mm_interconnect_0_onchip_memory2_0_s1_write),                  //                                           .write
		.onchip_memory2_0_s1_readdata                     (mm_interconnect_0_onchip_memory2_0_s1_readdata),               //                                           .readdata
		.onchip_memory2_0_s1_writedata                    (mm_interconnect_0_onchip_memory2_0_s1_writedata),              //                                           .writedata
		.onchip_memory2_0_s1_byteenable                   (mm_interconnect_0_onchip_memory2_0_s1_byteenable),             //                                           .byteenable
		.onchip_memory2_0_s1_chipselect                   (mm_interconnect_0_onchip_memory2_0_s1_chipselect),             //                                           .chipselect
		.onchip_memory2_0_s1_clken                        (mm_interconnect_0_onchip_memory2_0_s1_clken),                  //                                           .clken
		.out_scanner_s1_address                           (mm_interconnect_0_out_scanner_s1_address),                     //                             out_scanner_s1.address
		.out_scanner_s1_write                             (mm_interconnect_0_out_scanner_s1_write),                       //                                           .write
		.out_scanner_s1_readdata                          (mm_interconnect_0_out_scanner_s1_readdata),                    //                                           .readdata
		.out_scanner_s1_writedata                         (mm_interconnect_0_out_scanner_s1_writedata),                   //                                           .writedata
		.out_scanner_s1_chipselect                        (mm_interconnect_0_out_scanner_s1_chipselect),                  //                                           .chipselect
		.out_SPS_s1_address                               (mm_interconnect_0_out_sps_s1_address),                         //                                 out_SPS_s1.address
		.out_SPS_s1_write                                 (mm_interconnect_0_out_sps_s1_write),                           //                                           .write
		.out_SPS_s1_readdata                              (mm_interconnect_0_out_sps_s1_readdata),                        //                                           .readdata
		.out_SPS_s1_writedata                             (mm_interconnect_0_out_sps_s1_writedata),                       //                                           .writedata
		.out_SPS_s1_chipselect                            (mm_interconnect_0_out_sps_s1_chipselect),                      //                                           .chipselect
		.readyToTransfer_s1_address                       (mm_interconnect_0_readytotransfer_s1_address),                 //                         readyToTransfer_s1.address
		.readyToTransfer_s1_readdata                      (mm_interconnect_0_readytotransfer_s1_readdata)                 //                                           .readdata
	);

	nios2_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (nios2_qsys_0_d_irq_irq)          //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                             // reset_in0.reset
		.reset_in1      (nios2_qsys_0_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (clk_clk),                                    //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),             // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),         //          .reset_req
		.reset_req_in0  (1'b0),                                       // (terminated)
		.reset_req_in1  (1'b0),                                       // (terminated)
		.reset_in2      (1'b0),                                       // (terminated)
		.reset_req_in2  (1'b0),                                       // (terminated)
		.reset_in3      (1'b0),                                       // (terminated)
		.reset_req_in3  (1'b0),                                       // (terminated)
		.reset_in4      (1'b0),                                       // (terminated)
		.reset_req_in4  (1'b0),                                       // (terminated)
		.reset_in5      (1'b0),                                       // (terminated)
		.reset_req_in5  (1'b0),                                       // (terminated)
		.reset_in6      (1'b0),                                       // (terminated)
		.reset_req_in6  (1'b0),                                       // (terminated)
		.reset_in7      (1'b0),                                       // (terminated)
		.reset_req_in7  (1'b0),                                       // (terminated)
		.reset_in8      (1'b0),                                       // (terminated)
		.reset_req_in8  (1'b0),                                       // (terminated)
		.reset_in9      (1'b0),                                       // (terminated)
		.reset_req_in9  (1'b0),                                       // (terminated)
		.reset_in10     (1'b0),                                       // (terminated)
		.reset_req_in10 (1'b0),                                       // (terminated)
		.reset_in11     (1'b0),                                       // (terminated)
		.reset_req_in11 (1'b0),                                       // (terminated)
		.reset_in12     (1'b0),                                       // (terminated)
		.reset_req_in12 (1'b0),                                       // (terminated)
		.reset_in13     (1'b0),                                       // (terminated)
		.reset_req_in13 (1'b0),                                       // (terminated)
		.reset_in14     (1'b0),                                       // (terminated)
		.reset_req_in14 (1'b0),                                       // (terminated)
		.reset_in15     (1'b0),                                       // (terminated)
		.reset_req_in15 (1'b0)                                        // (terminated)
	);

endmodule
